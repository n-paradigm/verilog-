module password_save(
    input clk,
    input rst_n,
    input [3:0] key_value,    // 按键值
    input key_valid,          // 按键有效
    input [15:0] new_pwd,     // 新设置的密码（来自密码设置模块）
    input pwd_save,           // 密码保存信号（来自密码设置模块）
    output reg [15:0] input_pwd, // 输入的4位密码（每4位存1个数字，共16位）
    output   pwd_match,     // 密码匹配标志
    output reg [15:0] saved_pwd// 存储的密码
);



// 内部信号：记录输入的数字个数
reg [2:0] pwd_cnt=3'd0;
// 存储密码初始化与更新（新增：通过pwd_save信号触发更新）
always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        saved_pwd <= 16'h1111;
    end else if(pwd_save) begin
        // 密码更新：将新设置的密码保存
        saved_pwd <= new_pwd;
    end
end

// 密码输入逻辑（右入左移：输入1→0001，输入2→0012，输入3→0123，输入4→1234）
always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        input_pwd <= 16'h0000;
        pwd_cnt <= 3'd0;
    end else if(key_valid) begin
        case(key_value)
            4'd0,4'd1,4'd2,4'd3,4'd4,
            4'd5,4'd6,4'd7,4'd8,4'd9: begin // 0-9数字键
                if(pwd_cnt < 3'd4) begin
                    // 左移4位，新数字放在最低4位
                    input_pwd <= {input_pwd[11:0], key_value};
                    pwd_cnt <= pwd_cnt + 1'b1;
                end else begin
                    // 第4位数字：覆盖最左位
                    input_pwd <= {12'd0, key_value};
                    pwd_cnt <= 3'd1; // 重置计数，可重新输入
                end
            end
            4'b1101: begin // C键：清除密码
                input_pwd <= 16'h0000;
                pwd_cnt <= 3'd0;
            end
            4'b1011: begin // B键：退格
                if(pwd_cnt > 3'd0) begin
                    // 右移4位，最高4位置0
                    input_pwd <= {4'h0, input_pwd[15:4]};
                    pwd_cnt <= pwd_cnt - 1'b1;
                end else begin
                    input_pwd <= input_pwd; // 无数字可退格
                end
            end
            default: begin // 其他键不处理
                input_pwd <= input_pwd;
                pwd_cnt <= pwd_cnt;
            end
        endcase
    end
end


assign pwd_match = (input_pwd == saved_pwd) ? 1'b1 : 1'b0;
endmodule

/**
// 密码匹配判断（仅当输入4位密码后，按下确认键时判断）
always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        pwd_match <= 1'b0;
//    end else if(key_valid && key_value == 4'b1010) begin // A键：确认
	 end 
    else begin
		if(key_valid && key_value == 4'b1010)begin
			pwd_match <= (input_pwd == saved_pwd) ? 1'b1 : 1'b0;
		end
		else begin
			pwd_match <= 1'b0;
		end
	end
end


endmodule
**/